1
0 6 4 1 3 r h 2 B 44 H
3 2 0 0 1 r 26 30 38 40 44 47 48 49 52 53 57 h 27 B 32 B 40 B
7 0 3 0 0 r h 15 B 42 B
0 0 1 13 3 r 16 24 h 22 H 50 H
5 7 1 8 0 3 4 4 1 10 3 4 2 2 2 3 1 11 0 12 3 11 4 9 0 5 0 11 4 9 1 4 2 5 3 6 2 3
